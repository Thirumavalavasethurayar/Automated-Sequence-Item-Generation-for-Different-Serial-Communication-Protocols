`ifndef BASIC_IF__SV
`define BASIC_IF__SV

`include "basic_defines.svh"
interface basic_if (input bit clk, rst_n);

   logic                    data;
 
endinterface : basic_if

`endif //BASIC_IF__SV
