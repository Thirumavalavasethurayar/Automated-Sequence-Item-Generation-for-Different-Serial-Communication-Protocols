`ifndef BASIC_DEFINES__SVH
`define BASIC_DEFINES__SVH
 
`endif //BASIC_DEFINES__SVH
