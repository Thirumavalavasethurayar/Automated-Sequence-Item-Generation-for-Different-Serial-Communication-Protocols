`ifndef BASIC_PKG__SV
`define BASIC_PKG__SV
package basic_pkg;

  import uvm_pkg::*;
   `include "uvm_macros.svh"
   `include "basic_defines.svh"
   `include "basic_txn.svh"
   `include "basic_agent_cfg.svh"
   `include "basic_driver.svh"
   `include "basic_monitor.svh"
   `include "basic_agent.svh"

endpackage 
`endif //BASIC_PKG__SV
